`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Cal Poly 
// Engineer: Miguel Villa Floran
// 
// Create Date: 07/21/2024 11:49:15 AM
// Module Name: Arithmetic Logic Unit (ALU)
// Description: 
//////////////////////////////////////////////////////////////////////////////////

